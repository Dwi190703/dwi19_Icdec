magic
tech sky130A
magscale 1 2
timestamp 1729134742
<< nwell >>
rect -425 -1373 425 1373
<< pmos >>
rect -229 754 -29 1154
rect 29 754 229 1154
rect -229 118 -29 518
rect 29 118 229 518
rect -229 -518 -29 -118
rect 29 -518 229 -118
rect -229 -1154 -29 -754
rect 29 -1154 229 -754
<< pdiff >>
rect -287 1142 -229 1154
rect -287 766 -275 1142
rect -241 766 -229 1142
rect -287 754 -229 766
rect -29 1142 29 1154
rect -29 766 -17 1142
rect 17 766 29 1142
rect -29 754 29 766
rect 229 1142 287 1154
rect 229 766 241 1142
rect 275 766 287 1142
rect 229 754 287 766
rect -287 506 -229 518
rect -287 130 -275 506
rect -241 130 -229 506
rect -287 118 -229 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 229 506 287 518
rect 229 130 241 506
rect 275 130 287 506
rect 229 118 287 130
rect -287 -130 -229 -118
rect -287 -506 -275 -130
rect -241 -506 -229 -130
rect -287 -518 -229 -506
rect -29 -130 29 -118
rect -29 -506 -17 -130
rect 17 -506 29 -130
rect -29 -518 29 -506
rect 229 -130 287 -118
rect 229 -506 241 -130
rect 275 -506 287 -130
rect 229 -518 287 -506
rect -287 -766 -229 -754
rect -287 -1142 -275 -766
rect -241 -1142 -229 -766
rect -287 -1154 -229 -1142
rect -29 -766 29 -754
rect -29 -1142 -17 -766
rect 17 -1142 29 -766
rect -29 -1154 29 -1142
rect 229 -766 287 -754
rect 229 -1142 241 -766
rect 275 -1142 287 -766
rect 229 -1154 287 -1142
<< pdiffc >>
rect -275 766 -241 1142
rect -17 766 17 1142
rect 241 766 275 1142
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect -275 -506 -241 -130
rect -17 -506 17 -130
rect 241 -506 275 -130
rect -275 -1142 -241 -766
rect -17 -1142 17 -766
rect 241 -1142 275 -766
<< nsubdiff >>
rect -389 1303 -293 1337
rect 293 1303 389 1337
rect -389 1241 -355 1303
rect 355 1241 389 1303
rect -389 -1303 -355 -1241
rect 355 -1303 389 -1241
rect -389 -1337 -293 -1303
rect 293 -1337 389 -1303
<< nsubdiffcont >>
rect -293 1303 293 1337
rect -389 -1241 -355 1241
rect 355 -1241 389 1241
rect -293 -1337 293 -1303
<< poly >>
rect -229 1235 -29 1251
rect -229 1201 -213 1235
rect -45 1201 -29 1235
rect -229 1154 -29 1201
rect 29 1235 229 1251
rect 29 1201 45 1235
rect 213 1201 229 1235
rect 29 1154 229 1201
rect -229 707 -29 754
rect -229 673 -213 707
rect -45 673 -29 707
rect -229 657 -29 673
rect 29 707 229 754
rect 29 673 45 707
rect 213 673 229 707
rect 29 657 229 673
rect -229 599 -29 615
rect -229 565 -213 599
rect -45 565 -29 599
rect -229 518 -29 565
rect 29 599 229 615
rect 29 565 45 599
rect 213 565 229 599
rect 29 518 229 565
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect -229 -565 -29 -518
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect -229 -615 -29 -599
rect 29 -565 229 -518
rect 29 -599 45 -565
rect 213 -599 229 -565
rect 29 -615 229 -599
rect -229 -673 -29 -657
rect -229 -707 -213 -673
rect -45 -707 -29 -673
rect -229 -754 -29 -707
rect 29 -673 229 -657
rect 29 -707 45 -673
rect 213 -707 229 -673
rect 29 -754 229 -707
rect -229 -1201 -29 -1154
rect -229 -1235 -213 -1201
rect -45 -1235 -29 -1201
rect -229 -1251 -29 -1235
rect 29 -1201 229 -1154
rect 29 -1235 45 -1201
rect 213 -1235 229 -1201
rect 29 -1251 229 -1235
<< polycont >>
rect -213 1201 -45 1235
rect 45 1201 213 1235
rect -213 673 -45 707
rect 45 673 213 707
rect -213 565 -45 599
rect 45 565 213 599
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -599 -45 -565
rect 45 -599 213 -565
rect -213 -707 -45 -673
rect 45 -707 213 -673
rect -213 -1235 -45 -1201
rect 45 -1235 213 -1201
<< locali >>
rect -389 1303 -293 1337
rect 293 1303 389 1337
rect -389 1241 -355 1303
rect 355 1241 389 1303
rect -229 1201 -213 1235
rect -45 1201 -29 1235
rect 29 1201 45 1235
rect 213 1201 229 1235
rect -275 1142 -241 1158
rect -275 750 -241 766
rect -17 1142 17 1158
rect -17 750 17 766
rect 241 1142 275 1158
rect 241 750 275 766
rect -229 673 -213 707
rect -45 673 -29 707
rect 29 673 45 707
rect 213 673 229 707
rect -229 565 -213 599
rect -45 565 -29 599
rect 29 565 45 599
rect 213 565 229 599
rect -275 506 -241 522
rect -275 114 -241 130
rect -17 506 17 522
rect -17 114 17 130
rect 241 506 275 522
rect 241 114 275 130
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -130 -241 -114
rect -275 -522 -241 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 241 -130 275 -114
rect 241 -522 275 -506
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect 29 -599 45 -565
rect 213 -599 229 -565
rect -229 -707 -213 -673
rect -45 -707 -29 -673
rect 29 -707 45 -673
rect 213 -707 229 -673
rect -275 -766 -241 -750
rect -275 -1158 -241 -1142
rect -17 -766 17 -750
rect -17 -1158 17 -1142
rect 241 -766 275 -750
rect 241 -1158 275 -1142
rect -229 -1235 -213 -1201
rect -45 -1235 -29 -1201
rect 29 -1235 45 -1201
rect 213 -1235 229 -1201
rect -389 -1303 -355 -1241
rect 355 -1303 389 -1241
rect -389 -1337 -293 -1303
rect 293 -1337 389 -1303
<< viali >>
rect -213 1201 -45 1235
rect 45 1201 213 1235
rect -275 766 -241 1142
rect -17 766 17 1142
rect 241 766 275 1142
rect -213 673 -45 707
rect 45 673 213 707
rect -213 565 -45 599
rect 45 565 213 599
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -275 -506 -241 -130
rect -17 -506 17 -130
rect 241 -506 275 -130
rect -213 -599 -45 -565
rect 45 -599 213 -565
rect -213 -707 -45 -673
rect 45 -707 213 -673
rect -275 -1142 -241 -766
rect -17 -1142 17 -766
rect 241 -1142 275 -766
rect -213 -1235 -45 -1201
rect 45 -1235 213 -1201
<< metal1 >>
rect -225 1235 -33 1241
rect -225 1201 -213 1235
rect -45 1201 -33 1235
rect -225 1195 -33 1201
rect 33 1235 225 1241
rect 33 1201 45 1235
rect 213 1201 225 1235
rect 33 1195 225 1201
rect -281 1142 -235 1154
rect -281 766 -275 1142
rect -241 766 -235 1142
rect -281 754 -235 766
rect -23 1142 23 1154
rect -23 766 -17 1142
rect 17 766 23 1142
rect -23 754 23 766
rect 235 1142 281 1154
rect 235 766 241 1142
rect 275 766 281 1142
rect 235 754 281 766
rect -225 707 -33 713
rect -225 673 -213 707
rect -45 673 -33 707
rect -225 667 -33 673
rect 33 707 225 713
rect 33 673 45 707
rect 213 673 225 707
rect 33 667 225 673
rect -225 599 -33 605
rect -225 565 -213 599
rect -45 565 -33 599
rect -225 559 -33 565
rect 33 599 225 605
rect 33 565 45 599
rect 213 565 225 599
rect 33 559 225 565
rect -281 506 -235 518
rect -281 130 -275 506
rect -241 130 -235 506
rect -281 118 -235 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 235 506 281 518
rect 235 130 241 506
rect 275 130 281 506
rect 235 118 281 130
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect -281 -130 -235 -118
rect -281 -506 -275 -130
rect -241 -506 -235 -130
rect -281 -518 -235 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 235 -130 281 -118
rect 235 -506 241 -130
rect 275 -506 281 -130
rect 235 -518 281 -506
rect -225 -565 -33 -559
rect -225 -599 -213 -565
rect -45 -599 -33 -565
rect -225 -605 -33 -599
rect 33 -565 225 -559
rect 33 -599 45 -565
rect 213 -599 225 -565
rect 33 -605 225 -599
rect -225 -673 -33 -667
rect -225 -707 -213 -673
rect -45 -707 -33 -673
rect -225 -713 -33 -707
rect 33 -673 225 -667
rect 33 -707 45 -673
rect 213 -707 225 -673
rect 33 -713 225 -707
rect -281 -766 -235 -754
rect -281 -1142 -275 -766
rect -241 -1142 -235 -766
rect -281 -1154 -235 -1142
rect -23 -766 23 -754
rect -23 -1142 -17 -766
rect 17 -1142 23 -766
rect -23 -1154 23 -1142
rect 235 -766 281 -754
rect 235 -1142 241 -766
rect 275 -1142 281 -766
rect 235 -1154 281 -1142
rect -225 -1201 -33 -1195
rect -225 -1235 -213 -1201
rect -45 -1235 -33 -1201
rect -225 -1241 -33 -1235
rect 33 -1201 225 -1195
rect 33 -1235 45 -1201
rect 213 -1235 225 -1201
rect 33 -1241 225 -1235
<< properties >>
string FIXED_BBOX -372 -1320 372 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
