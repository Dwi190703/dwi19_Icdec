magic
tech sky130A
magscale 1 2
timestamp 1729344248
<< nwell >>
rect -335 -914 810 746
rect -335 -915 90 -914
rect 181 -915 810 -914
rect -335 -1922 810 -915
<< pdiff >>
rect 184 -1233 230 -1221
<< nsubdiff >>
rect -299 676 -239 710
rect 714 676 774 710
rect -299 650 -265 676
rect 740 650 774 676
rect -299 -1852 -265 -1826
rect 740 -1852 774 -1826
rect -299 -1886 -239 -1852
rect 714 -1886 774 -1852
<< nsubdiffcont >>
rect -239 676 714 710
rect -299 -1826 -265 650
rect 740 -1826 774 650
rect -239 -1886 714 -1852
<< poly >>
rect 6 66 36 113
rect -59 50 36 66
rect -59 16 -43 50
rect -9 16 36 50
rect -59 0 36 16
rect 410 67 440 111
rect 410 51 506 67
rect 410 17 456 51
rect 490 17 506 51
rect 410 1 506 17
rect 5 -441 35 -397
rect -58 -457 35 -441
rect -58 -491 -42 -457
rect -8 -491 35 -457
rect -58 -507 35 -491
rect 409 -441 439 -399
rect 409 -457 503 -441
rect 409 -491 453 -457
rect 487 -491 503 -457
rect -58 -630 32 -614
rect 93 -617 191 -503
rect 251 -617 348 -504
rect 409 -507 503 -491
rect -58 -664 -42 -630
rect -8 -664 32 -630
rect -58 -680 32 -664
rect 2 -724 32 -680
rect 406 -630 502 -614
rect 406 -664 452 -630
rect 486 -664 502 -630
rect 406 -680 502 -664
rect 406 -730 436 -680
rect -62 -1137 33 -1121
rect -62 -1171 -46 -1137
rect -12 -1171 33 -1137
rect -62 -1187 33 -1171
rect 3 -1245 33 -1187
rect 407 -1137 503 -1121
rect 407 -1171 453 -1137
rect 487 -1171 503 -1137
rect 407 -1187 503 -1171
rect 407 -1243 437 -1187
<< polycont >>
rect -43 16 -9 50
rect 456 17 490 51
rect -42 -491 -8 -457
rect 453 -491 487 -457
rect -42 -664 -8 -630
rect 452 -664 486 -630
rect -46 -1171 -12 -1137
rect 453 -1171 487 -1137
<< locali >>
rect -299 676 -239 710
rect 714 676 774 710
rect -299 650 -265 676
rect 740 650 774 676
rect -59 16 -43 50
rect -9 16 7 50
rect 440 17 456 51
rect 490 17 506 51
rect -58 -491 -42 -457
rect -8 -491 8 -457
rect 437 -491 453 -457
rect 487 -491 503 -457
rect -58 -664 -42 -630
rect -8 -664 8 -630
rect 436 -664 452 -630
rect 486 -664 502 -630
rect -62 -1171 -46 -1137
rect -12 -1171 4 -1137
rect 437 -1171 453 -1137
rect 487 -1171 503 -1137
rect -299 -1852 -265 -1826
rect 740 -1852 774 -1826
rect -299 -1886 -239 -1852
rect 714 -1886 774 -1852
<< viali >>
rect 33 676 303 710
rect 33 675 303 676
rect -43 16 -9 50
rect 456 17 490 51
rect -42 -491 -8 -457
rect 453 -491 487 -457
rect -42 -664 -8 -630
rect 452 -664 486 -630
rect -46 -1171 -12 -1137
rect 453 -1171 487 -1137
<< metal1 >>
rect 21 710 315 716
rect 21 675 33 710
rect 303 675 315 710
rect 21 669 315 675
rect 455 586 510 592
rect 0 531 455 586
rect 0 300 55 531
rect 455 525 510 531
rect -50 100 89 300
rect 186 112 196 288
rect 248 112 258 288
rect 355 100 400 300
rect 452 100 496 300
rect -50 56 -1 100
rect -55 50 3 56
rect -55 16 -43 50
rect -9 16 3 50
rect -55 10 3 16
rect 122 -19 166 19
rect 258 11 268 63
rect 336 11 346 63
rect 450 57 495 100
rect 444 51 502 57
rect 444 17 456 51
rect 490 17 502 51
rect 444 11 502 17
rect 450 10 495 11
rect 121 -63 328 -19
rect 99 -169 109 -117
rect 177 -169 187 -117
rect 284 -126 328 -63
rect -50 -219 89 -206
rect 356 -219 495 -205
rect -50 -395 -49 -219
rect 3 -395 89 -219
rect 185 -395 195 -219
rect 247 -395 257 -219
rect 356 -395 441 -219
rect 493 -395 503 -219
rect -50 -406 89 -395
rect 356 -405 495 -395
rect -46 -451 -1 -406
rect 445 -451 492 -405
rect -54 -457 4 -451
rect -54 -491 -42 -457
rect -8 -491 4 -457
rect -54 -497 4 -491
rect 441 -457 499 -451
rect 441 -491 453 -457
rect 487 -491 499 -457
rect 441 -497 499 -491
rect -46 -498 -1 -497
rect -50 -624 -5 -623
rect -54 -630 4 -624
rect -54 -664 -42 -630
rect -8 -664 4 -630
rect -54 -670 4 -664
rect 440 -630 498 -624
rect 440 -664 452 -630
rect 486 -664 498 -630
rect 440 -670 498 -664
rect -50 -715 -5 -670
rect 448 -714 482 -670
rect -51 -726 90 -715
rect -62 -902 -52 -726
rect 0 -902 90 -726
rect 190 -726 242 -715
rect 354 -726 489 -714
rect 190 -727 194 -726
rect -51 -915 90 -902
rect 181 -902 194 -727
rect 246 -902 256 -726
rect 354 -902 439 -726
rect 491 -902 501 -726
rect 181 -915 242 -902
rect 354 -915 489 -902
rect 96 -1003 106 -951
rect 174 -1003 184 -951
rect 265 -1033 326 -973
rect 113 -1094 326 -1033
rect -58 -1137 0 -1131
rect -58 -1171 -46 -1137
rect -12 -1171 0 -1137
rect 113 -1158 174 -1094
rect -58 -1177 0 -1171
rect -46 -1221 -4 -1177
rect 255 -1184 265 -1132
rect 333 -1184 343 -1132
rect 441 -1137 499 -1131
rect 441 -1171 453 -1137
rect 487 -1171 499 -1137
rect 441 -1177 499 -1171
rect 448 -1221 489 -1177
rect -52 -1422 86 -1221
rect 197 -1233 249 -1221
rect 183 -1409 193 -1233
rect 245 -1409 249 -1233
rect 197 -1421 249 -1409
rect 349 -1233 489 -1221
rect 349 -1409 440 -1233
rect 492 -1409 502 -1233
rect 349 -1421 489 -1409
rect -9 -1646 54 -1422
rect 448 -1646 529 -1636
rect -9 -1709 455 -1646
rect 518 -1709 529 -1646
rect 448 -1716 529 -1709
<< via1 >>
rect 455 531 510 586
rect 196 112 248 288
rect 400 100 452 300
rect 268 11 336 63
rect 109 -169 177 -117
rect -49 -395 3 -219
rect 195 -395 247 -219
rect 441 -395 493 -219
rect -52 -902 0 -726
rect 194 -902 246 -726
rect 439 -902 491 -726
rect 106 -1003 174 -951
rect 265 -1184 333 -1132
rect 193 -1409 245 -1233
rect 440 -1409 492 -1233
rect 455 -1709 518 -1646
<< metal2 >>
rect 453 589 513 598
rect 449 531 453 586
rect 513 531 516 586
rect 453 520 513 529
rect -52 424 452 476
rect -52 -209 0 424
rect 400 300 452 424
rect 196 288 252 298
rect 196 102 252 112
rect 400 90 452 100
rect 268 63 336 73
rect 268 1 336 11
rect 283 -27 328 1
rect 121 -72 328 -27
rect 121 -107 166 -72
rect 109 -117 177 -107
rect 109 -179 177 -169
rect -52 -219 3 -209
rect -52 -395 -49 -219
rect -52 -405 3 -395
rect 193 -219 249 -209
rect 193 -405 249 -395
rect 439 -219 495 -209
rect 439 -405 495 -395
rect -52 -726 0 -405
rect -52 -1548 0 -902
rect 191 -726 247 -716
rect 191 -912 247 -902
rect 438 -726 494 -716
rect 438 -912 494 -902
rect 106 -951 174 -941
rect 106 -1013 174 -1003
rect 113 -1039 174 -1013
rect 113 -1095 326 -1039
rect 265 -1122 326 -1095
rect 265 -1132 333 -1122
rect 265 -1194 333 -1184
rect 445 -1223 497 -1219
rect 191 -1233 247 -1223
rect 191 -1419 247 -1409
rect 440 -1233 497 -1223
rect 492 -1409 497 -1233
rect 440 -1419 497 -1409
rect 445 -1548 497 -1419
rect -52 -1600 497 -1548
rect 448 -1646 525 -1636
rect 448 -1709 455 -1646
rect 518 -1709 525 -1646
rect 448 -1715 525 -1709
<< via2 >>
rect 453 586 513 589
rect 453 531 455 586
rect 455 531 510 586
rect 510 531 513 586
rect 453 529 513 531
rect 196 112 248 288
rect 248 112 252 288
rect 193 -395 195 -219
rect 195 -395 247 -219
rect 247 -395 249 -219
rect 439 -395 441 -219
rect 441 -395 493 -219
rect 493 -395 495 -219
rect 191 -902 194 -726
rect 194 -902 246 -726
rect 246 -902 247 -726
rect 438 -902 439 -726
rect 439 -902 491 -726
rect 491 -902 494 -726
rect 191 -1409 193 -1233
rect 193 -1409 245 -1233
rect 245 -1409 247 -1233
rect 458 -1706 514 -1650
<< metal3 >>
rect 448 589 518 594
rect 448 529 453 589
rect 513 529 518 589
rect 448 524 518 529
rect 186 288 262 293
rect 186 146 196 288
rect 174 112 196 146
rect 252 146 262 288
rect 453 242 513 524
rect 252 112 267 146
rect 174 -219 267 112
rect 452 -214 514 242
rect 429 -219 514 -214
rect 174 -235 193 -219
rect 181 -395 193 -235
rect 249 -236 266 -219
rect 249 -395 259 -236
rect 181 -400 259 -395
rect 429 -395 439 -219
rect 495 -232 514 -219
rect 495 -395 516 -232
rect 429 -400 516 -395
rect 181 -726 258 -400
rect 453 -489 516 -400
rect 453 -513 517 -489
rect 454 -641 517 -513
rect 454 -721 519 -641
rect 181 -902 191 -726
rect 247 -902 258 -726
rect 181 -1233 258 -902
rect 428 -726 519 -721
rect 428 -902 438 -726
rect 494 -871 519 -726
rect 494 -902 520 -871
rect 428 -907 520 -902
rect 455 -1233 520 -907
rect 181 -1409 191 -1233
rect 247 -1409 258 -1233
rect 181 -1415 258 -1409
rect 448 -1645 522 -1233
rect 453 -1650 519 -1645
rect 453 -1706 458 -1650
rect 514 -1706 519 -1650
rect 453 -1711 519 -1706
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729240092
transform 1 0 20 0 1 -307
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729240092
transform 1 0 18 0 1 -1321
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729240092
transform 1 0 422 0 1 -1321
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729240092
transform 1 0 17 0 1 -814
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729240092
transform 1 0 421 0 1 -814
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729240092
transform 1 0 424 0 1 -307
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729240092
transform 1 0 425 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729240092
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729238916
transform 1 0 220 0 1 -1321
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729238916
transform 1 0 223 0 1 200
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_2
timestamp 1729238916
transform 1 0 222 0 1 -307
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_3
timestamp 1729238916
transform 1 0 219 0 1 -814
box -223 -200 223 200
<< labels >>
flabel viali 153 695 153 695 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal2 77 445 77 445 0 FreeSans 800 0 0 0 D6
port 1 nsew
flabel metal1 156 -9 156 -9 0 FreeSans 800 0 0 0 VIP
port 2 nsew
flabel metal2 149 -82 149 -82 0 FreeSans 800 0 0 0 VIN
port 3 nsew
flabel metal3 218 -148 218 -148 0 FreeSans 800 0 0 0 D5
port 4 nsew
flabel metal3 485 418 485 418 0 FreeSans 800 0 0 0 OUT
port 5 nsew
<< end >>
