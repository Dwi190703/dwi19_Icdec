magic
tech sky130A
magscale 1 2
timestamp 1729218920
<< error_p >>
rect -194 18 194 236
<< nwell >>
rect -194 18 194 618
rect -194 -618 194 -18
<< pmos >>
rect -100 118 100 518
rect -100 -518 100 -118
<< pdiff >>
rect -158 506 -100 518
rect -158 130 -146 506
rect -112 130 -100 506
rect -158 118 -100 130
rect 100 506 158 518
rect 100 130 112 506
rect 146 130 158 506
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -506 -146 -130
rect -112 -506 -100 -130
rect -158 -518 -100 -506
rect 100 -130 158 -118
rect 100 -506 112 -130
rect 146 -506 158 -130
rect 100 -518 158 -506
<< pdiffc >>
rect -146 130 -112 506
rect 112 130 146 506
rect -146 -506 -112 -130
rect 112 -506 146 -130
<< poly >>
rect -100 599 100 615
rect -100 565 -84 599
rect 84 565 100 599
rect -100 518 100 565
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -565 100 -518
rect -100 -599 -84 -565
rect 84 -599 100 -565
rect -100 -615 100 -599
<< polycont >>
rect -84 565 84 599
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -599 84 -565
<< locali >>
rect -100 565 -84 599
rect 84 565 100 599
rect -146 506 -112 522
rect -146 114 -112 130
rect 112 506 146 522
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -522 -112 -506
rect 112 -130 146 -114
rect 112 -522 146 -506
rect -100 -599 -84 -565
rect 84 -599 100 -565
<< viali >>
rect -84 565 84 599
rect -146 130 -112 506
rect 112 130 146 506
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -506 -112 -130
rect 112 -506 146 -130
rect -84 -599 84 -565
<< metal1 >>
rect -96 599 96 605
rect -96 565 -84 599
rect 84 565 96 599
rect -96 559 96 565
rect -152 506 -106 518
rect -152 130 -146 506
rect -112 130 -106 506
rect -152 118 -106 130
rect 106 506 152 518
rect 106 130 112 506
rect 146 130 152 506
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -506 -146 -130
rect -112 -506 -106 -130
rect -152 -518 -106 -506
rect 106 -130 152 -118
rect 106 -506 112 -130
rect 146 -506 152 -130
rect 106 -518 152 -506
rect -96 -565 96 -559
rect -96 -599 -84 -565
rect 84 -599 96 -565
rect -96 -605 96 -599
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
