magic
tech sky130A
magscale 1 2
timestamp 1729422980
<< metal1 >>
rect 2079 3339 2131 3345
rect 2079 3281 2131 3287
rect -890 3105 -838 3111
rect -890 3047 -838 3053
rect -884 2704 -850 3047
rect 1575 2791 1618 2796
rect 90 2757 1618 2791
rect 2088 2789 2122 3281
rect 2263 3222 3466 3258
rect 2263 2789 2299 3222
rect 2765 3052 2771 3104
rect 2823 3052 2829 3104
rect 2780 2926 2814 3052
rect -880 2589 -852 2704
rect 90 1965 124 2757
rect 1575 2561 1618 2757
rect 1540 2551 1618 2561
rect 1332 2518 1618 2551
rect 1332 2517 1567 2518
rect -669 1931 124 1965
rect 1767 2088 2130 2122
rect 1653 1942 1659 1943
rect 1585 1922 1659 1942
rect 1331 1892 1659 1922
rect 1331 1890 1591 1892
rect 1653 1891 1659 1892
rect 1711 1891 1717 1943
rect 590 1680 625 1761
rect 590 1673 628 1680
rect 591 1623 628 1673
rect 1296 1636 1350 1638
rect 592 1565 627 1623
rect 1286 1584 1296 1636
rect 1352 1584 1362 1636
rect 592 1530 774 1565
rect 739 1402 774 1530
rect -24 1297 352 1300
rect -77 1266 352 1297
rect 1296 1280 1350 1584
rect -77 1264 25 1266
rect -77 1263 -1 1264
rect -836 918 -174 953
rect -77 -277 -43 1263
rect 1767 -277 1801 2088
rect 2052 -172 2104 -166
rect 3430 -178 3466 3222
rect 2104 -218 3468 -178
rect 3430 -220 3466 -218
rect 2052 -230 2104 -224
rect -77 -311 1801 -277
<< via1 >>
rect 2079 3287 2131 3339
rect -890 3053 -838 3105
rect 2771 3052 2823 3104
rect 1659 1891 1711 1943
rect 1296 1584 1352 1636
rect 2052 -224 2104 -172
<< metal2 >>
rect 3528 3342 3593 3352
rect 2073 3287 2079 3339
rect 2131 3287 3528 3339
rect 3528 3268 3593 3278
rect -896 3053 -890 3105
rect -838 3104 -832 3105
rect 2771 3104 2823 3110
rect -838 3054 2771 3104
rect -838 3053 -832 3054
rect 2823 3054 2825 3104
rect 2771 3046 2823 3052
rect 1655 2920 1716 2930
rect 1655 2809 1716 2859
rect 1660 1949 1710 2809
rect 1659 1943 1711 1949
rect -797 1842 -223 1887
rect 1659 1885 1711 1891
rect 1296 1638 1352 1646
rect 1296 1636 1392 1638
rect 892 1213 926 1589
rect 1352 1626 1392 1636
rect 1352 1586 1662 1626
rect 1296 1574 1352 1584
rect 1622 -178 1662 1586
rect 2046 -178 2052 -172
rect 1622 -218 2052 -178
rect 2046 -224 2052 -218
rect 2104 -224 2110 -172
<< via2 >>
rect 3528 3278 3593 3342
rect 1655 2859 1716 2920
<< metal3 >>
rect 3518 3342 3603 3347
rect 3518 3278 3528 3342
rect 3593 3278 3603 3342
rect 3518 3273 3603 3278
rect 1645 2920 1726 2925
rect -19 2859 1655 2920
rect 1716 2859 1726 2920
rect -19 1830 42 2859
rect 1645 2854 1726 2859
rect -643 1769 42 1830
rect -934 -461 -870 520
rect 3528 -461 3592 3273
rect -934 -525 3592 -461
use nmos2  nmos2_0
timestamp 1729346615
transform 1 0 360 0 1 2186
box -208 -442 1155 528
use nmoscs  nmoscs_0
timestamp 1729224578
transform 1 0 -794 0 1 92
box 794 -92 2654 1349
use pmos2  pmos2_0
timestamp 1729344248
transform 1 0 -1125 0 1 1914
box -335 -1922 810 746
use pmoscs  pmoscs_0
timestamp 1729359038
transform 1 0 2129 0 1 837
box -249 -833 916 2158
<< labels >>
flabel metal3 12 2874 12 2874 0 FreeSans 1600 0 0 0 out
port 1 nsew
flabel metal2 910 1498 910 1498 0 FreeSans 1600 0 0 0 rs
port 2 nsew
flabel metal1 -254 940 -254 940 0 FreeSans 1600 0 0 0 vip
port 3 nsew
flabel metal2 -262 1860 -262 1860 0 FreeSans 1600 0 0 0 vin
port 4 nsew
flabel metal1 612 1602 612 1602 0 FreeSans 1600 0 0 0 gnd
port 5 nsew
flabel metal2 -528 3076 -528 3076 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
<< end >>
