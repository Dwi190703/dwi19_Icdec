magic
tech sky130A
magscale 1 2
timestamp 1729218920
<< nmos >>
rect -100 47 100 447
rect -100 -447 100 -47
<< ndiff >>
rect -158 435 -100 447
rect -158 59 -146 435
rect -112 59 -100 435
rect -158 47 -100 59
rect 100 435 158 447
rect 100 59 112 435
rect 146 59 158 435
rect 100 47 158 59
rect -158 -59 -100 -47
rect -158 -435 -146 -59
rect -112 -435 -100 -59
rect -158 -447 -100 -435
rect 100 -59 158 -47
rect 100 -435 112 -59
rect 146 -435 158 -59
rect 100 -447 158 -435
<< ndiffc >>
rect -146 59 -112 435
rect 112 59 146 435
rect -146 -435 -112 -59
rect 112 -435 146 -59
<< poly >>
rect -100 447 100 473
rect -100 21 100 47
rect -100 -47 100 -21
rect -100 -473 100 -447
<< locali >>
rect -146 435 -112 451
rect -146 43 -112 59
rect 112 435 146 451
rect 112 43 146 59
rect -146 -59 -112 -43
rect -146 -451 -112 -435
rect 112 -59 146 -43
rect 112 -451 146 -435
<< viali >>
rect -146 59 -112 435
rect 112 59 146 435
rect -146 -435 -112 -59
rect 112 -435 146 -59
<< metal1 >>
rect -152 435 -106 447
rect -152 59 -146 435
rect -112 59 -106 435
rect -152 47 -106 59
rect 106 435 152 447
rect 106 59 112 435
rect 146 59 152 435
rect 106 47 152 59
rect -152 -59 -106 -47
rect -152 -435 -146 -59
rect -112 -435 -106 -59
rect -152 -447 -106 -435
rect 106 -59 152 -47
rect 106 -435 112 -59
rect 146 -435 152 -59
rect 106 -447 152 -435
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
