magic
tech sky130A
magscale 1 2
timestamp 1729224578
<< psubdiff >>
rect 905 1309 965 1343
rect 2309 1309 2369 1343
rect 905 1283 939 1309
rect 2335 1283 2369 1309
rect 905 -52 939 -26
rect 2335 -52 2369 -26
rect 905 -86 965 -52
rect 2309 -86 2369 -52
<< psubdiffcont >>
rect 965 1309 2309 1343
rect 905 -26 939 1283
rect 2335 -26 2369 1283
rect 965 -86 2309 -52
<< poly >>
rect 1496 1173 1757 1212
rect 1321 586 1932 648
rect 1505 24 1766 63
<< locali >>
rect 905 1309 965 1343
rect 2309 1309 2369 1343
rect 905 1283 939 1309
rect 905 -52 939 -26
rect 2335 1283 2369 1309
rect 2335 -52 2369 -26
rect 905 -86 965 -52
rect 2309 -86 2369 -52
<< viali >>
rect 1533 1309 1567 1343
rect 1686 -86 1720 -52
<< metal1 >>
rect 1521 1343 1579 1349
rect 1521 1309 1533 1343
rect 1567 1309 1579 1343
rect 1521 1303 1579 1309
rect 1074 1127 1109 1217
rect 1159 1127 1312 1130
rect 1074 1116 1312 1127
rect 1533 1121 1567 1303
rect 2128 1206 2178 1210
rect 2124 1187 2178 1206
rect 2124 1168 2181 1187
rect 1940 1124 2093 1129
rect 2152 1124 2181 1168
rect 1075 763 1312 1116
rect 1075 748 1315 763
rect 1159 746 1315 748
rect 1269 703 1315 746
rect 1269 701 1316 703
rect 1269 655 1355 701
rect 1533 638 1567 760
rect 1667 748 1677 1124
rect 1729 748 1739 1124
rect 1925 748 1935 1124
rect 1987 1116 2181 1124
rect 1987 748 2178 1116
rect 1940 745 2178 748
rect 1533 604 1720 638
rect 1159 489 1312 490
rect 1075 486 1312 489
rect 1075 110 1263 486
rect 1315 110 1325 486
rect 1514 110 1524 486
rect 1576 110 1586 486
rect 1686 474 1720 604
rect 1891 536 1978 570
rect 1941 490 1978 536
rect 1939 486 2092 490
rect 1075 20 1112 110
rect 1159 106 1312 110
rect 1686 -46 1720 130
rect 1939 107 2179 486
rect 1939 106 2093 107
rect 2047 68 2093 106
rect 2046 10 2110 68
rect 1674 -52 1732 -46
rect 1674 -86 1686 -52
rect 1720 -86 1732 -52
rect 1674 -92 1732 -86
<< via1 >>
rect 1677 748 1729 1124
rect 1935 748 1987 1124
rect 1263 110 1315 486
rect 1524 110 1576 486
<< metal2 >>
rect 1677 1124 1729 1134
rect 1677 738 1729 748
rect 1933 1124 1989 1134
rect 1933 738 1989 748
rect 1686 637 1720 738
rect 1534 603 1720 637
rect 1534 598 1568 603
rect 1533 496 1567 598
rect 1261 486 1317 496
rect 1261 100 1317 110
rect 1524 486 1576 496
rect 1524 100 1576 110
<< via2 >>
rect 1933 748 1935 1124
rect 1935 748 1987 1124
rect 1987 748 1989 1124
rect 1261 110 1263 486
rect 1263 110 1315 486
rect 1315 110 1317 486
<< metal3 >>
rect 1923 1124 1999 1129
rect 1923 748 1933 1124
rect 1989 748 1999 1124
rect 1923 743 1999 748
rect 1935 651 1995 743
rect 1254 590 1996 651
rect 1254 491 1315 590
rect 1935 589 1995 590
rect 1251 486 1327 491
rect 1251 110 1261 486
rect 1317 110 1327 486
rect 1251 105 1327 110
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_0
timestamp 1729218920
transform 1 0 1421 0 1 936
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_1
timestamp 1729218920
transform 1 0 1421 0 1 298
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_2
timestamp 1729218920
transform 1 0 1832 0 1 298
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_3
timestamp 1729218920
transform 1 0 1832 0 1 936
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_L2VWCK  sky130_fd_pr__nfet_01v8_L2VWCK_0
timestamp 1729224578
transform 1 0 2117 0 1 267
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_LG94FM  sky130_fd_pr__nfet_01v8_LG94FM_0
timestamp 1729224578
transform 1 0 2117 0 1 967
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_LG94FM  sky130_fd_pr__nfet_01v8_LG94FM_1
timestamp 1729224578
transform 1 0 1136 0 1 967
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_SCJFGL  sky130_fd_pr__nfet_01v8_SCJFGL_0
timestamp 1729224578
transform 1 0 1136 0 1 267
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_TCR5KT  sky130_fd_pr__nfet_01v8_TCR5KT_1
timestamp 1729218920
transform 1 0 2653 0 1 755
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_TCR5KT  sky130_fd_pr__nfet_01v8_TCR5KT_2
timestamp 1729218920
transform 1 0 2392 0 1 532
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_TCR5KT  sky130_fd_pr__nfet_01v8_TCR5KT_3
timestamp 1729218920
transform 1 0 794 0 1 410
box 0 0 1 1
<< labels >>
flabel metal1 1287 712 1287 712 0 FreeSans 1600 0 0 0 d3
port 0 nsew
flabel metal2 1702 679 1702 679 0 FreeSans 1600 0 0 0 rs
port 1 nsew
flabel metal3 1968 660 1968 660 0 FreeSans 1600 0 0 0 d4
port 2 nsew
flabel metal1 1699 -25 1699 -25 0 FreeSans 1600 0 0 0 gnd
port 3 nsew
<< end >>
